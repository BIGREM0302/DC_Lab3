module AudPlayer();


endmodule